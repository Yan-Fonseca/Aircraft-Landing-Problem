module main
import file_manager {read_data}

fn main() {
	read_data("/home/iamthemage/Documentos/Aircraft-Landing-Problem/instances/airland1.txt")
}
