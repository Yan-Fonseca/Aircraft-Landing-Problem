module constructive

