module main
import file_manager {read_data}

fn main() {
	read_data("/home/yan/inteligencia_computacional/ALP/instances/airland1.txt")
}
