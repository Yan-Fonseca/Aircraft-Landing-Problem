module filemanager
import os
import models

pub fn read_data(path string) Problem {
	mut counter := 0
	lines := read_lines(path)
	for line in lines { 
		// realizar a leitura dos arquivos
	}
}